// define enumerated types for packet payload size
`define SMALL 0
`define MEDIUM 1
`define LARGE 2

module generator();

reg [0:7] uid; 								// Unique id field to identify the packet
reg [7:0] len;
reg [7:0] Da, rand_port;
reg [7:0] Sa;
reg [0:7] pkt [0:258]; 				// Maximum packet size (259 8-bit Bytes)
reg [0:7] parity;

integer payload_size;					// Control field for the payload size
integer parity_type;					// Control field for the parity type

initial
	uid = 0;


task randomize();
	begin
		uid = uid + 1;
		parity_type = {$random}%2;		// 0 and 1 are selected randomly
		rand_port = {$random}%4;			// 0, 1, 2, and 3 are selected randomly
		Da = $root.tbench_top.test.env.mem[rand_port];
		Sa = $random;

		if ( $root.tbench_top.test.randomize_payload_size == 1 ) begin
			payload_size = {$random}%3;		// 0, 1, and 2 are selected randomly
			if ( payload_size == `SMALL )
				len = {$random}%10;					// payload between 0-9 bytes
			else if ( payload_size == `MEDIUM )
				len = 10 + {$random}%10;		// payload between 10-19 bytes
			else if ( payload_size == `LARGE )
				len = 20 + {$random}%10;		// payload between 20-29 bytes
			else
				len = 30 + {$random}%10;		// payload between 30-39 bytes
			end

		else
			len = $root.tbench_top.test.env.size_of_payload;

		if ( parity_type == 0 )
			parity = 8'b0;
		else
			parity = 8'b1;

	end
endtask


task packing();
	integer i;
	begin
		pkt[0] = Da;		// port it should be going to
		pkt[1] = Sa;		// port it's coming from
		pkt[2] = len;		// length of generated bytes (payload length)
		$display("[PACKING] pkt[0] is Da %b %d, Sa %b %d, len %b %d ", pkt[0], Da, Sa, Sa, len, len);

		for ( i=0; i<len+3; i=i+1 )
			pkt[i+3] = $random;

		pkt[3] = uid;
		pkt[i+3] = parity ^ parity_cal(0);

	end
endtask


function [0:7] parity_cal(input_dummy);
	integer i;
	reg [0:7] result;
	begin
		result = 8'hFF;
		for ( i=0; i<len+4; i=i+1 )
			begin
				result = result ^ pkt[i];
			end
		parity_cal=result;

	end
endfunction


endmodule
