`ifndef TESTBENCH_SV
`define TESTBENCH_SV

program testbench(intf i_intf);

  initial
  begin
    $display("******************* Start of testcase ****************");
  end

endprogram

`endif
