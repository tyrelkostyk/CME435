program testbench (
// interface and ports here...   
);

// testbench code here...

initial begin
  $display("Running test_sanity...");
  // ...
  // ...
end 

endprogram
