program testbench( intf i_intf );

initial begin
	$display("*************** Start of testbench ***************");
end

final
	$display("*************** End of testbench ***************");


endprogram
